VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO low_swing_tx
  CLASS CORE ;
  ORIGIN -0.8 -0.5 ;
  FOREIGN low_swing_tx 0.8 0.5 ;
  SIZE 33.08 BY 2.205 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vss
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.04 0.5 33.6 0.83 ;
        RECT 27.57 0.5 27.66 1.245 ;
        RECT 22.08 0.5 22.17 1.245 ;
        RECT 16.14 0.5 16.23 1.245 ;
        RECT 14.46 0.5 14.55 1.245 ;
        RECT 12.78 0.5 12.87 1.245 ;
        RECT 6.94 0.5 7.03 1.245 ;
        RECT 5.26 0.5 5.35 1.245 ;
        RECT 3.58 0.5 3.67 1.245 ;
        RECT 1.98 0.5 2.07 1.245 ;
    END
  END vss
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2 1.555 1.685 1.645 ;
        RECT 1.2 1.555 1.29 1.89 ;
    END
  END i
  PIN vdd
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.04 2.3 33.6 2.63 ;
        RECT 27.98 1.775 28.07 2.63 ;
        RECT 27.16 1.775 27.25 2.63 ;
        RECT 26.34 1.775 26.43 2.63 ;
        RECT 25.52 1.775 25.61 2.63 ;
        RECT 24.7 1.775 24.79 2.63 ;
        RECT 23.88 1.775 23.97 2.63 ;
        RECT 22.9 1.775 22.99 2.63 ;
        RECT 22.08 1.775 22.17 2.63 ;
        RECT 21.18 1.775 21.27 2.63 ;
        RECT 19.5 1.775 19.59 2.63 ;
        RECT 17.82 1.775 17.91 2.63 ;
        RECT 16.14 1.775 16.23 2.63 ;
        RECT 14.46 1.775 14.55 2.63 ;
        RECT 12.78 1.775 12.87 2.63 ;
        RECT 11.98 1.775 12.07 2.63 ;
        RECT 10.3 1.775 10.39 2.63 ;
        RECT 8.62 1.775 8.71 2.63 ;
        RECT 6.94 1.775 7.03 2.63 ;
        RECT 5.26 1.775 5.35 2.63 ;
        RECT 3.58 1.775 3.67 2.63 ;
        RECT 2.8 1.775 2.89 2.63 ;
        RECT 1.98 1.775 2.07 2.63 ;
    END
  END vdd
  PIN c
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 32.67 1.555 32.76 1.945 ;
        RECT 29.39 1.555 32.76 1.645 ;
        RECT 31.85 1.555 31.94 1.945 ;
        RECT 31.03 1.555 31.12 1.945 ;
        RECT 30.21 1.1 30.69 1.19 ;
        RECT 30.21 0.955 30.3 1.945 ;
        RECT 27.98 0.955 30.3 1.045 ;
        RECT 29.39 1.555 29.48 1.945 ;
        RECT 27.98 0.955 28.07 1.245 ;
    END
  END c
  OBS
    LAYER M1 ;
      RECT 28.455 2.055 33.17 2.145 ;
      RECT 33.08 1.775 33.17 2.145 ;
      RECT 32.26 1.775 32.35 2.145 ;
      RECT 31.44 1.775 31.53 2.145 ;
      RECT 30.62 1.775 30.71 2.145 ;
      RECT 29.8 1.775 29.89 2.145 ;
      RECT 28.98 1.555 29.07 2.145 ;
      RECT 28.455 1.555 28.545 2.145 ;
      RECT 27.57 1.555 27.66 1.945 ;
      RECT 26.75 1.555 26.84 1.945 ;
      RECT 25.93 1.555 26.02 1.945 ;
      RECT 25.11 1.555 25.2 1.945 ;
      RECT 24.29 1.555 24.38 1.945 ;
      RECT 24.29 1.555 28.545 1.645 ;
      RECT 22.49 1.075 22.58 1.945 ;
      RECT 22.49 1.355 29.315 1.445 ;
      RECT 23.21 1.55 23.39 1.65 ;
      RECT 23.21 1.555 23.785 1.645 ;
      RECT 20.34 1.555 20.43 1.945 ;
      RECT 18.66 1.555 18.75 1.945 ;
      RECT 16.98 1.075 17.07 1.945 ;
      RECT 15.3 1.555 15.39 1.945 ;
      RECT 13.62 1.555 13.71 1.945 ;
      RECT 13.62 1.555 21.685 1.645 ;
      RECT 13.62 1.355 17.07 1.445 ;
      RECT 15.3 1.075 15.39 1.445 ;
      RECT 13.62 1.075 13.71 1.445 ;
      RECT 11.14 1.555 11.23 1.945 ;
      RECT 9.46 1.555 9.55 1.945 ;
      RECT 7.78 1.075 7.87 1.945 ;
      RECT 6.1 1.555 6.19 1.945 ;
      RECT 4.42 1.555 4.51 1.945 ;
      RECT 4.42 1.555 12.385 1.645 ;
      RECT 4.42 1.355 7.87 1.445 ;
      RECT 6.1 1.075 6.19 1.445 ;
      RECT 4.42 1.075 4.51 1.445 ;
      RECT 2.39 1.075 2.48 1.945 ;
      RECT 2.39 1.455 3.185 1.545 ;
      RECT 10.715 1.05 11.19 1.15 ;
    LAYER M2 ;
      RECT 23.25 1.35 23.35 1.69 ;
      RECT 11.05 1.35 23.35 1.45 ;
      RECT 11.05 1.01 11.15 1.45 ;
    LAYER VIA1 ;
      RECT 23.25 1.55 23.35 1.65 ;
      RECT 11.05 1.05 11.15 1.15 ;
  END
END low_swing_tx

END LIBRARY

* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d0 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_CDNS_733622483252
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nch_CDNS_733622483254
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pch_CDNS_733622483251
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nch_CDNS_733622483250
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_CDNS_733622483252
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pch_CDNS_733622483253
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT low_swing_tx vss vdd c i
** N=9 EP=4 IP=45 FDC=57
M0 3 i vss vss nch L=6e-08 W=1.2e-07 $X=2200 $Y=1100 $D=6
M1 6 3 vss vss nch L=4.9e-07 W=1.2e-07 $X=3800 $Y=1100 $D=6
M2 vss 3 6 vss nch L=4.9e-07 W=1.2e-07 $X=4640 $Y=1100 $D=6
M3 6 3 vss vss nch L=4.9e-07 W=1.2e-07 $X=5480 $Y=1100 $D=6
M4 vss 3 6 vss nch L=4.9e-07 W=1.2e-07 $X=6320 $Y=1100 $D=6
M5 6 3 vss vss nch L=4.9e-07 W=1.2e-07 $X=7160 $Y=1100 $D=6
M6 7 6 vss vss nch L=4.9e-07 W=1.2e-07 $X=13000 $Y=1100 $D=6
M7 vss 6 7 vss nch L=4.9e-07 W=1.2e-07 $X=13840 $Y=1100 $D=6
M8 7 6 vss vss nch L=4.9e-07 W=1.2e-07 $X=14680 $Y=1100 $D=6
M9 vss 6 7 vss nch L=4.9e-07 W=1.2e-07 $X=15520 $Y=1100 $D=6
M10 7 6 vss vss nch L=4.9e-07 W=1.2e-07 $X=16360 $Y=1100 $D=6
M11 4 7 vss vss nch L=6e-08 W=1.2e-07 $X=22300 $Y=1100 $D=6
M12 c 3 vss vss nch L=6e-08 W=1.2e-07 $X=27790 $Y=1100 $D=6
M13 3 i vdd vdd pch L=6e-08 W=1.2e-07 $X=2200 $Y=1800 $D=101
M14 vdd i 3 vdd pch L=6e-08 W=1.2e-07 $X=2610 $Y=1800 $D=101
M15 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=3800 $Y=1800 $D=101
M16 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 $X=4640 $Y=1800 $D=101
M17 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=5480 $Y=1800 $D=101
M18 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 $X=6320 $Y=1800 $D=101
M19 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=7160 $Y=1800 $D=101
M20 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 $X=8000 $Y=1800 $D=101
M21 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=8840 $Y=1800 $D=101
M22 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 $X=9680 $Y=1800 $D=101
M23 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=10520 $Y=1800 $D=101
M24 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 $X=11360 $Y=1800 $D=101
M25 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=13000 $Y=1800 $D=101
M26 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 $X=13840 $Y=1800 $D=101
M27 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=14680 $Y=1800 $D=101
M28 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 $X=15520 $Y=1800 $D=101
M29 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=16360 $Y=1800 $D=101
M30 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 $X=17200 $Y=1800 $D=101
M31 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=18040 $Y=1800 $D=101
M32 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 $X=18880 $Y=1800 $D=101
M33 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 $X=19720 $Y=1800 $D=101
M34 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 $X=20560 $Y=1800 $D=101
M35 4 7 vdd vdd pch L=6e-08 W=1.2e-07 $X=22300 $Y=1800 $D=101
M36 vdd 7 4 vdd pch L=6e-08 W=1.2e-07 $X=22710 $Y=1800 $D=101
M37 8 3 vdd vdd pch L=6e-08 W=1.2e-07 $X=24100 $Y=1800 $D=101
M38 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 $X=24510 $Y=1800 $D=101
M39 8 3 vdd vdd pch L=6e-08 W=1.2e-07 $X=24920 $Y=1800 $D=101
M40 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 $X=25330 $Y=1800 $D=101
M41 8 3 vdd vdd pch L=6e-08 W=1.2e-07 $X=25740 $Y=1800 $D=101
M42 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 $X=26150 $Y=1800 $D=101
M43 8 3 vdd vdd pch L=6e-08 W=1.2e-07 $X=26560 $Y=1800 $D=101
M44 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 $X=26970 $Y=1800 $D=101
M45 8 3 vdd vdd pch L=6e-08 W=1.2e-07 $X=27380 $Y=1800 $D=101
M46 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 $X=27790 $Y=1800 $D=101
M47 c 4 8 vdd pch L=6e-08 W=1.2e-07 $X=29200 $Y=1800 $D=101
M48 8 4 c vdd pch L=6e-08 W=1.2e-07 $X=29610 $Y=1800 $D=101
M49 c 4 8 vdd pch L=6e-08 W=1.2e-07 $X=30020 $Y=1800 $D=101
M50 8 4 c vdd pch L=6e-08 W=1.2e-07 $X=30430 $Y=1800 $D=101
M51 c 4 8 vdd pch L=6e-08 W=1.2e-07 $X=30840 $Y=1800 $D=101
M52 8 4 c vdd pch L=6e-08 W=1.2e-07 $X=31250 $Y=1800 $D=101
M53 c 4 8 vdd pch L=6e-08 W=1.2e-07 $X=31660 $Y=1800 $D=101
M54 8 4 c vdd pch L=6e-08 W=1.2e-07 $X=32070 $Y=1800 $D=101
M55 c 4 8 vdd pch L=6e-08 W=1.2e-07 $X=32480 $Y=1800 $D=101
M56 8 4 c vdd pch L=6e-08 W=1.2e-07 $X=32890 $Y=1800 $D=101
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d0 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_CDNS_733622498682
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nch_CDNS_733622498684
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pch_CDNS_733622498681
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nch_CDNS_733622498680
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_CDNS_733622498682
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pch_CDNS_733622498683
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT low_swing_tx vss vdd c i
** N=9 EP=4 IP=37 FDC=57
M0 3 i vss vss nch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=3.45e-14 PD=8e-07 PS=8e-07 NRD=2.39583 NRS=2.39583 sa=2.5e-07 sb=2.5e-07 sca=11.7338 scb=0.0125229 scc=0.000446911 $X=2200 $Y=1100 $D=6
M1 6 3 vss vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=3.61e-06 sca=11.3401 scb=0.012522 scc=0.000446911 $X=3800 $Y=1100 $D=6
M2 vss 3 6 vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.09e-06 sb=2.77e-06 sca=11.3048 scb=0.012522 scc=0.000446911 $X=4640 $Y=1100 $D=6
M3 6 3 vss vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.93e-06 sb=1.93e-06 sca=11.2861 scb=0.012522 scc=0.000446911 $X=5480 $Y=1100 $D=6
M4 vss 3 6 vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.77e-06 sb=1.09e-06 sca=11.2813 scb=0.012522 scc=0.000446911 $X=6320 $Y=1100 $D=6
M5 6 3 vss vss nch L=4.9e-07 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=3.61e-06 sb=2.5e-07 sca=11.2813 scb=0.012522 scc=0.000446911 $X=7160 $Y=1100 $D=6
M6 7 6 vss vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=3.61e-06 sca=11.2813 scb=0.012522 scc=0.000446911 $X=13000 $Y=1100 $D=6
M7 vss 6 7 vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.09e-06 sb=2.77e-06 sca=11.2813 scb=0.012522 scc=0.000446911 $X=13840 $Y=1100 $D=6
M8 7 6 vss vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.93e-06 sb=1.93e-06 sca=11.2813 scb=0.012522 scc=0.000446911 $X=14680 $Y=1100 $D=6
M9 vss 6 7 vss nch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.77e-06 sb=1.09e-06 sca=11.2813 scb=0.012522 scc=0.000446911 $X=15520 $Y=1100 $D=6
M10 7 6 vss vss nch L=4.9e-07 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=3.61e-06 sb=2.5e-07 sca=11.2813 scb=0.012522 scc=0.000446911 $X=16360 $Y=1100 $D=6
M11 4 7 vss vss nch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=3.45e-14 PD=8e-07 PS=8e-07 NRD=2.39583 NRS=2.39583 sa=2.5e-07 sb=2.5e-07 sca=11.2875 scb=0.012522 scc=0.000446911 $X=22300 $Y=1100 $D=6
M12 c 3 vss vss nch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=3.45e-14 PD=8e-07 PS=8e-07 NRD=2.39583 NRS=2.39583 sa=2.5e-07 sb=2.5e-07 sca=11.2875 scb=0.012522 scc=0.000446911 $X=27790 $Y=1100 $D=6
M13 3 i vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=6.6e-07 sca=9.87288 scb=0.0102876 scc=0.000317496 $X=2200 $Y=1800 $D=101
M14 vdd i 3 vdd pch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=6.6e-07 sb=2.5e-07 sca=9.67909 scb=0.0102868 scc=0.000317496 $X=2610 $Y=1800 $D=101
M15 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=7.81e-06 sca=9.47606 scb=0.0102867 scc=0.000317496 $X=3800 $Y=1800 $D=101
M16 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.09e-06 sb=6.97e-06 sca=9.44069 scb=0.0102867 scc=0.000317496 $X=4640 $Y=1800 $D=101
M17 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.93e-06 sb=6.13e-06 sca=9.42188 scb=0.0102867 scc=0.000317496 $X=5480 $Y=1800 $D=101
M18 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.77e-06 sb=5.29e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=6320 $Y=1800 $D=101
M19 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.61e-06 sb=4.45e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=7160 $Y=1800 $D=101
M20 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=4.45e-06 sb=3.61e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=8000 $Y=1800 $D=101
M21 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=5.29e-06 sb=2.77e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=8840 $Y=1800 $D=101
M22 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.13e-06 sb=1.93e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=9680 $Y=1800 $D=101
M23 6 3 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.97e-06 sb=1.09e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=10520 $Y=1800 $D=101
M24 vdd 3 6 vdd pch L=4.9e-07 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=7.81e-06 sb=2.5e-07 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=11360 $Y=1800 $D=101
M25 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=7.81e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=13000 $Y=1800 $D=101
M26 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.09e-06 sb=6.97e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=13840 $Y=1800 $D=101
M27 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.93e-06 sb=6.13e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=14680 $Y=1800 $D=101
M28 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.77e-06 sb=5.29e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=15520 $Y=1800 $D=101
M29 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.61e-06 sb=4.45e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=16360 $Y=1800 $D=101
M30 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=4.45e-06 sb=3.61e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=17200 $Y=1800 $D=101
M31 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=5.29e-06 sb=2.77e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=18040 $Y=1800 $D=101
M32 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.13e-06 sb=1.93e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=18880 $Y=1800 $D=101
M33 7 6 vdd vdd pch L=4.9e-07 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.97e-06 sb=1.09e-06 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=19720 $Y=1800 $D=101
M34 vdd 6 7 vdd pch L=4.9e-07 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=7.81e-06 sb=2.5e-07 sca=9.41698 scb=0.0102867 scc=0.000317496 $X=20560 $Y=1800 $D=101
M35 4 7 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=6.6e-07 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=22300 $Y=1800 $D=101
M36 vdd 7 4 vdd pch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=6.6e-07 sb=2.5e-07 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=22710 $Y=1800 $D=101
M37 8 3 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=3.94e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=24100 $Y=1800 $D=101
M38 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.6e-07 sb=3.53e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=24510 $Y=1800 $D=101
M39 8 3 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.07e-06 sb=3.12e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=24920 $Y=1800 $D=101
M40 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.48e-06 sb=2.71e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=25330 $Y=1800 $D=101
M41 8 3 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.89e-06 sb=2.3e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=25740 $Y=1800 $D=101
M42 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.3e-06 sb=1.89e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=26150 $Y=1800 $D=101
M43 8 3 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.71e-06 sb=1.48e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=26560 $Y=1800 $D=101
M44 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.12e-06 sb=1.07e-06 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=26970 $Y=1800 $D=101
M45 8 3 vdd vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.53e-06 sb=6.6e-07 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=27380 $Y=1800 $D=101
M46 vdd 3 8 vdd pch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=3.94e-06 sb=2.5e-07 sca=9.42317 scb=0.0102867 scc=0.000317496 $X=27790 $Y=1800 $D=101
M47 c 4 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=3.45e-14 PD=5e-07 PS=8e-07 NRD=1.61458 NRS=2.39583 sa=2.5e-07 sb=3.94e-06 sca=9.42989 scb=0.0102867 scc=0.000317496 $X=29200 $Y=1800 $D=101
M48 8 4 c vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=6.6e-07 sb=3.53e-06 sca=9.43927 scb=0.0102867 scc=0.000317496 $X=29610 $Y=1800 $D=101
M49 c 4 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.07e-06 sb=3.12e-06 sca=9.45182 scb=0.0102867 scc=0.000317496 $X=30020 $Y=1800 $D=101
M50 8 4 c vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.48e-06 sb=2.71e-06 sca=9.46914 scb=0.0102867 scc=0.000317496 $X=30430 $Y=1800 $D=101
M51 c 4 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=1.89e-06 sb=2.3e-06 sca=9.49403 scb=0.0102867 scc=0.000317496 $X=30840 $Y=1800 $D=101
M52 8 4 c vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.3e-06 sb=1.89e-06 sca=9.53159 scb=0.0102867 scc=0.000317496 $X=31250 $Y=1800 $D=101
M53 c 4 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=2.71e-06 sb=1.48e-06 sca=9.59218 scb=0.0102867 scc=0.000317496 $X=31660 $Y=1800 $D=101
M54 8 4 c vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.12e-06 sb=1.07e-06 sca=9.69935 scb=0.0102868 scc=0.000317496 $X=32070 $Y=1800 $D=101
M55 c 4 8 vdd pch L=6e-08 W=1.2e-07 AD=2.325e-14 AS=2.325e-14 PD=5e-07 PS=5e-07 NRD=1.61458 NRS=1.61458 sa=3.53e-06 sb=6.6e-07 sca=9.91669 scb=0.0102883 scc=0.000317496 $X=32480 $Y=1800 $D=101
M56 8 4 c vdd pch L=6e-08 W=1.2e-07 AD=3.45e-14 AS=2.325e-14 PD=8e-07 PS=5e-07 NRD=2.39583 NRS=1.61458 sa=3.94e-06 sb=2.5e-07 sca=10.4698 scb=0.0103525 scc=0.0003175 $X=32890 $Y=1800 $D=101
.ENDS
***************************************

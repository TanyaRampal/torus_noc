** Generated for: hspiceD
** Generated on: Dec  5 22:06:23 2024
** Design library name: ece720t7
** Design cell name: torus_xbar_1b
** Design view name: schematic


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/CMC/tsmc_65nm/CRN65GP/TN65CMSP018K3_V1.0C/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt

** Library name: ece720t7
** Cell name: torus_xbar_1b
** View name: schematic
.subckt torus_xbar_1b eo n2s ni p2e p2s pi so vss w2e w2s wi
m4 ni n2s so vss nch l=60e-9 w=200e-9 m=1 nf=1 sd=200e-9 ad=35e-15 as=35e-15 pd=750e-9 ps=750e-9 nrd=500e-3 nrs=500e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m3 wi w2s so vss nch l=60e-9 w=200e-9 m=1 nf=1 sd=200e-9 ad=35e-15 as=35e-15 pd=750e-9 ps=750e-9 nrd=500e-3 nrs=500e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m2 pi p2s so vss nch l=60e-9 w=200e-9 m=1 nf=1 sd=200e-9 ad=35e-15 as=35e-15 pd=750e-9 ps=750e-9 nrd=500e-3 nrs=500e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m1 pi p2e eo vss nch l=60e-9 w=200e-9 m=1 nf=1 sd=200e-9 ad=35e-15 as=35e-15 pd=750e-9 ps=750e-9 nrd=500e-3 nrs=500e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m0 wi w2e eo vss nch l=60e-9 w=200e-9 m=1 nf=1 sd=200e-9 ad=35e-15 as=35e-15 pd=750e-9 ps=750e-9 nrd=500e-3 nrs=500e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends torus_xbar_1b
** End of subcircuit definition.
.END

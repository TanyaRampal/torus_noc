`timescale 1ns/1ps


module low_swing_rx (
    input wire i,
    output wire o
);

assign o = i;

endmodule

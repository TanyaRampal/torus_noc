`timescale 1ns/1ps

module low_swing_tx (
    input wire i,
    output wire c
);

assign c = i;

endmodule

